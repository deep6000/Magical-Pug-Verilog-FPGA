// VGA_Subsystem.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module VGA_Subsystem (
		input  wire       clk_clk,         //     clk.clk
		output wire [7:0] digit_0_digit_0, // digit_0.digit_0
		output wire [7:0] digit_1_digit_1, // digit_1.digit_1
		output wire [7:0] digit_2_digit_2, // digit_2.digit_2
		input  wire [3:0] keys_keys,       //    keys.keys
		input  wire       reset_reset_n,   //   reset.reset_n
		output wire [7:0] score_score,     //   score.score
		input  wire       switch_switch,   //  switch.switch
		output wire       vga_CLK,         //     vga.CLK
		output wire       vga_HS,          //        .HS
		output wire       vga_VS,          //        .VS
		output wire       vga_BLANK,       //        .BLANK
		output wire       vga_SYNC,        //        .SYNC
		output wire [7:0] vga_R,           //        .R
		output wire [7:0] vga_G,           //        .G
		output wire [7:0] vga_B            //        .B
	);

	wire         vga_fifo_avalon_dc_buffer_source_valid;                        // vga_fifo:stream_out_valid -> vga_controller:valid
	wire  [29:0] vga_fifo_avalon_dc_buffer_source_data;                         // vga_fifo:stream_out_data -> vga_controller:data
	wire         vga_fifo_avalon_dc_buffer_source_ready;                        // vga_controller:ready -> vga_fifo:stream_out_ready
	wire         vga_fifo_avalon_dc_buffer_source_startofpacket;                // vga_fifo:stream_out_startofpacket -> vga_controller:startofpacket
	wire         vga_fifo_avalon_dc_buffer_source_endofpacket;                  // vga_fifo:stream_out_endofpacket -> vga_controller:endofpacket
	wire         rgb_resampler_avalon_rgb_source_valid;                         // rgb_resampler:stream_out_valid -> vga_fifo:stream_in_valid
	wire  [29:0] rgb_resampler_avalon_rgb_source_data;                          // rgb_resampler:stream_out_data -> vga_fifo:stream_in_data
	wire         rgb_resampler_avalon_rgb_source_ready;                         // vga_fifo:stream_in_ready -> rgb_resampler:stream_out_ready
	wire         rgb_resampler_avalon_rgb_source_startofpacket;                 // rgb_resampler:stream_out_startofpacket -> vga_fifo:stream_in_startofpacket
	wire         rgb_resampler_avalon_rgb_source_endofpacket;                   // rgb_resampler:stream_out_endofpacket -> vga_fifo:stream_in_endofpacket
	wire         video_pll_0_vga_clk_clk;                                       // video_pll_0:vga_clk_clk -> [rst_controller_001:clk, rst_controller_002:clk, vga_controller:clk, vga_fifo:clk_stream_out]
	wire         magical_pug_generator_0_avalon_streaming_source_valid;         // magical_pug_generator_0:valid -> avalon_st_adapter:in_0_valid
	wire  [23:0] magical_pug_generator_0_avalon_streaming_source_data;          // magical_pug_generator_0:data -> avalon_st_adapter:in_0_data
	wire         magical_pug_generator_0_avalon_streaming_source_ready;         // avalon_st_adapter:in_0_ready -> magical_pug_generator_0:ready
	wire         magical_pug_generator_0_avalon_streaming_source_startofpacket; // magical_pug_generator_0:startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         magical_pug_generator_0_avalon_streaming_source_endofpacket;   // magical_pug_generator_0:endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire   [1:0] magical_pug_generator_0_avalon_streaming_source_empty;         // magical_pug_generator_0:empty -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                                 // avalon_st_adapter:out_0_valid -> rgb_resampler:stream_in_valid
	wire  [23:0] avalon_st_adapter_out_0_data;                                  // avalon_st_adapter:out_0_data -> rgb_resampler:stream_in_data
	wire         avalon_st_adapter_out_0_ready;                                 // rgb_resampler:stream_in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                         // avalon_st_adapter:out_0_startofpacket -> rgb_resampler:stream_in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                           // avalon_st_adapter:out_0_endofpacket -> rgb_resampler:stream_in_endofpacket
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, magical_pug_generator_0:reset, rgb_resampler:reset, vga_fifo:reset_stream_in]
	wire         rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> vga_controller:reset
	wire         rst_controller_002_reset_out_reset;                            // rst_controller_002:reset_out -> vga_fifo:reset_stream_out
	wire         video_pll_0_reset_source_reset;                                // video_pll_0:reset_source_reset -> rst_controller_002:reset_in0

	magical_pug_generator #(
		.DW     (23),
		.WW     (10),
		.HW     (9),
		.WIDTH  (640),
		.HEIGHT (480)
	) magical_pug_generator_0 (
		.clk           (clk_clk),                                                       //                   clock.clk
		.reset         (rst_controller_reset_out_reset),                                //                   reset.reset
		.ready         (magical_pug_generator_0_avalon_streaming_source_ready),         // avalon_streaming_source.ready
		.data          (magical_pug_generator_0_avalon_streaming_source_data),          //                        .data
		.startofpacket (magical_pug_generator_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.endofpacket   (magical_pug_generator_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.empty         (magical_pug_generator_0_avalon_streaming_source_empty),         //                        .empty
		.valid         (magical_pug_generator_0_avalon_streaming_source_valid),         //                        .valid
		.keys          (keys_keys),                                                     //                    keys.keys
		.score         (score_score),                                                   //                   score.score
		.switch        (switch_switch),                                                 //                  switch.switch
		.digit_0       (digit_0_digit_0),                                               //                 Digit_0.digit_0
		.digit_1       (digit_1_digit_1),                                               //                 Digit_1.digit_1
		.digit_2       (digit_2_digit_2)                                                //                 Digit_2.digit_2
	);

	VGA_Subsystem_rgb_resampler rgb_resampler (
		.clk                      (clk_clk),                                       //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                //             reset.reset
		.stream_in_startofpacket  (avalon_st_adapter_out_0_startofpacket),         //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (avalon_st_adapter_out_0_endofpacket),           //                  .endofpacket
		.stream_in_valid          (avalon_st_adapter_out_0_valid),                 //                  .valid
		.stream_in_ready          (avalon_st_adapter_out_0_ready),                 //                  .ready
		.stream_in_data           (avalon_st_adapter_out_0_data),                  //                  .data
		.slave_read               (),                                              //  avalon_rgb_slave.read
		.slave_readdata           (),                                              //                  .readdata
		.stream_out_ready         (rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	VGA_Subsystem_vga_controller vga_controller (
		.clk           (video_pll_0_vga_clk_clk),                        //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),             //              reset.reset
		.data          (vga_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (vga_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (vga_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (vga_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (vga_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                                        // external_interface.export
		.VGA_HS        (vga_HS),                                         //                   .export
		.VGA_VS        (vga_VS),                                         //                   .export
		.VGA_BLANK     (vga_BLANK),                                      //                   .export
		.VGA_SYNC      (vga_SYNC),                                       //                   .export
		.VGA_R         (vga_R),                                          //                   .export
		.VGA_G         (vga_G),                                          //                   .export
		.VGA_B         (vga_B)                                           //                   .export
	);

	VGA_Subsystem_vga_fifo vga_fifo (
		.clk_stream_in            (clk_clk),                                        //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                 //         reset_stream_in.reset
		.clk_stream_out           (video_pll_0_vga_clk_clk),                        //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),             //        reset_stream_out.reset
		.stream_in_ready          (rgb_resampler_avalon_rgb_source_ready),          //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (rgb_resampler_avalon_rgb_source_startofpacket),  //                        .startofpacket
		.stream_in_endofpacket    (rgb_resampler_avalon_rgb_source_endofpacket),    //                        .endofpacket
		.stream_in_valid          (rgb_resampler_avalon_rgb_source_valid),          //                        .valid
		.stream_in_data           (rgb_resampler_avalon_rgb_source_data),           //                        .data
		.stream_out_ready         (vga_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (vga_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (vga_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (vga_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (vga_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	VGA_Subsystem_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clk_clk),                        //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),                 //    ref_reset.reset
		.vga_clk_clk        (video_pll_0_vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (video_pll_0_reset_source_reset)  // reset_source.reset
	);

	VGA_Subsystem_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                                // in_rst_0.reset
		.in_0_data           (magical_pug_generator_0_avalon_streaming_source_data),          //     in_0.data
		.in_0_valid          (magical_pug_generator_0_avalon_streaming_source_valid),         //         .valid
		.in_0_ready          (magical_pug_generator_0_avalon_streaming_source_ready),         //         .ready
		.in_0_startofpacket  (magical_pug_generator_0_avalon_streaming_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (magical_pug_generator_0_avalon_streaming_source_endofpacket),   //         .endofpacket
		.in_0_empty          (magical_pug_generator_0_avalon_streaming_source_empty),         //         .empty
		.out_0_data          (avalon_st_adapter_out_0_data),                                  //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                                 //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                                 //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),                         //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)                            //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (video_pll_0_vga_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (video_pll_0_reset_source_reset),     // reset_in0.reset
		.clk            (video_pll_0_vga_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
